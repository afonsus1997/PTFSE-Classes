

module controller(
    input clock,
    input reset,
    input start,
    output init,
    output running,
    output toggle,
    output finish,
    output bist_end
    
);

//code here


endmodule // controller